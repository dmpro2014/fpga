library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package constants is
end;

package body constants is
	constant INSTRUCTION_ADDRESS_WIDTH = 16;
	constant WORD_WIDTH;
	end;
