library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity control_unit is
    Port ( instruction_in : in  STD_LOGIC_VECTOR (15 downto 0));
end control_unit;

architecture Behavioral of control_unit is

begin


end Behavioral;